LIBRARY IEEE;
USE IEEE.STD_Logic_1164.ALL;

ENTITY NAND_GATE IS
    PORT (
        A : IN STD_LOGIC;
        B : IN STD_LOGIC;
        Y : OUT STD_LOGIC
    );
END NAND_GATE;

ARCHITECTURE behavioural OF NAND_GATE IS
BEGIN

    Y <= A NAND B;
END behavioural;